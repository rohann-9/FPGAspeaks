`timescale 1ns / 1ps
module mux16x1_tb();
reg [15:0]d;
reg [3:0]s;
wire y;
mux16x1 DUT(d,s,y);
initial
begin
d=16'b1011010110001010;
s[3]=0;s[2]=0;s[1]=0;s[0]=0;#5
s[3]=0;s[2]=0;s[1]=0;s[0]=1;#5
s[3]=0;s[2]=0;s[1]=1;s[0]=0;#5
s[3]=0;s[2]=0;s[1]=1;s[0]=1;#5
s[3]=0;s[2]=1;s[1]=0;s[0]=0;#5
s[3]=0;s[2]=1;s[1]=0;s[0]=1;#5
s[3]=0;s[2]=1;s[1]=1;s[0]=0;#5
s[3]=0;s[2]=1;s[1]=1;s[0]=1;#5
s[3]=1;s[2]=0;s[1]=0;s[0]=0;#5
s[3]=1;s[2]=0;s[1]=0;s[0]=1;#5
s[3]=1;s[2]=0;s[1]=1;s[0]=0;#5
s[3]=1;s[2]=0;s[1]=1;s[0]=1;#5
s[3]=1;s[2]=1;s[1]=0;s[0]=0;#5
s[3]=1;s[2]=1;s[1]=0;s[0]=1;#5
s[3]=1;s[2]=1;s[1]=1;s[0]=0;#5
s[3]=1;s[2]=1;s[1]=1;s[0]=1;#5
$finish;
end
endmodule
