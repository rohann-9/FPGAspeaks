`timescale 1ns / 1ps
module q9_tb();
reg a,b,c,d;
wire f2;
q9 DUT(a,b,c,d,f2);
initial
begin
a=0;b=0;c=0;d=0;#10
a=0;b=0;c=0;d=1;#10
a=0;b=0;c=1;d=0;#10
a=0;b=0;c=1;d=1;#10
a=0;b=1;c=0;d=0;#10
a=0;b=1;c=0;d=1;#10
a=0;b=1;c=1;d=0;#10
a=0;b=1;c=1;d=1;#10
a=1;b=0;c=0;d=0;#10
a=1;b=0;c=0;d=1;#10
a=1;b=0;c=1;d=0;#10
a=1;b=0;c=1;d=1;#10
a=1;b=1;c=0;d=0;#10
a=1;b=1;c=0;d=1;#10
a=1;b=1;c=1;d=0;#10
a=1;b=1;c=1;d=1;#10
$finish;
end
endmodule
